***Phase_detector***
Vcdl 2 0 Pulse (5 0 5 0 0 10 20)
Vin 1 0 Pulse (5 0 0 0 0 10 20)
Vdd 3 0 DC 5

.model pmod pmos level=54 version=4.7 
.model nmod nmos level=54 version=4.7 

M1 4 1 3 3 pmod W = 20u  L = 1u 
M4 6 2 3 3 pmod W = 20u  L = 1u 
M7 5 4 1 1 pmod W = 20u  L = 1u 
M9 7 6 2 2 pmod W = 20u  L = 1u 
M11 10 5 1 1 pmod W = 20u  L = 1u 
M13 11 7 2 2 pmod W = 20u  L = 1u 

M2 4 1 8 8 nmod W = 10u L = 1u 
M5 6 2 9 9 nmod W = 10u L = 1u 
M3 8 2 0 0 nmod W = 10u L = 1u 
M6 9 1 0 0 nmod W = 10u L = 1u 
M8 5 4 0 0 nmod W = 10u L = 1u 
M10 7 6 0 0 nmod W = 10u L = 1u 
M12 10 5 0 0 nmod W = 10u L = 1u 
M14 11 7 0 0 nmod W = 10u L = 1u 

.tran 0.1 40
.control
run
plot V(1) title "IN"
plot V(2) title "VHDL"
plot V(10) title "Up"
plot V(11) title "Down"
.endc
.end
